module mux4_1_tb();

   //Step1 : Write down the variables required for testbench		
								
   //Step2 : Instantiate the Design 

   //Step3 : Declare a task to initialize inputs of DUT to 0 

   //Step4 : Declare  tasks with arguments for driving stimulus to DUT 

   //Step5 : Call the tasks from procedural process 

   //Step6 : Use $monitor task to display inputs and outputs

   //Step7 : Use $finish task to terminate the simulation at 100ns

   
endmodule

